// DE1_SOC_NIOS_2.v

// Generated using ACDS version 15.0 145

`timescale 1 ps / 1 ps
module DE1_SOC_NIOS_2 (
		input  wire        clk_clk,                           //                         clk.clk
		output wire        clock_23m_clk,                     //                   clock_23m.clk
		output wire        clock_6400k_clk,                   //                 clock_6400k.clk
		output wire        i2c_rst,                           //                         i2c.rst
		inout  wire        i2c_sda,                           //                            .sda
		inout  wire        i2c_sclk,                          //                            .sclk
		output wire [12:0] new_sdram_controller_0_wire_addr,  // new_sdram_controller_0_wire.addr
		output wire [1:0]  new_sdram_controller_0_wire_ba,    //                            .ba
		output wire        new_sdram_controller_0_wire_cas_n, //                            .cas_n
		output wire        new_sdram_controller_0_wire_cke,   //                            .cke
		output wire        new_sdram_controller_0_wire_cs_n,  //                            .cs_n
		inout  wire [15:0] new_sdram_controller_0_wire_dq,    //                            .dq
		output wire [1:0]  new_sdram_controller_0_wire_dqm,   //                            .dqm
		output wire        new_sdram_controller_0_wire_ras_n, //                            .ras_n
		output wire        new_sdram_controller_0_wire_we_n,  //                            .we_n
		input  wire        pixel_read_clk,                    //                       pixel.read_clk
		input  wire        pixel_ready,                       //                            .ready
		output wire        pixel_valid,                       //                            .valid
		output wire [15:0] pixel_readdata,                    //                            .readdata
		input  wire        pixel_frame_sync,                  //                            .frame_sync
		input  wire        reset_reset_n,                     //                       reset.reset_n
		output wire        sd_sd_cs,                          //                          sd.sd_cs
		output wire        sd_sd_clk,                         //                            .sd_clk
		output wire        sd_sd_di,                          //                            .sd_di
		input  wire        sd_sd_do,                          //                            .sd_do
		output wire        sdram_clk_clk                      //                   sdram_clk.clk
	);

	wire         pll_outclk0_clk;                                           // pll:outclk_0 -> [SPI_AVALON_SD_0:clk, cpu:clk, framebuffer_sdram_0:clk, i2c_AVALON_0:clk, irq_mapper:clk, jtag_uart:clk, mm_interconnect_0:pll_outclk0_clk, new_sdram_controller_0:clk, onchip_memory2:clk, rst_controller:clk]
	wire         framebuffer_sdram_0_avalon_master_chipselect;              // framebuffer_sdram_0:m0_chipselect -> mm_interconnect_0:framebuffer_sdram_0_avalon_master_chipselect
	wire         framebuffer_sdram_0_avalon_master_waitrequest;             // mm_interconnect_0:framebuffer_sdram_0_avalon_master_waitrequest -> framebuffer_sdram_0:m0_waitrequest
	wire  [15:0] framebuffer_sdram_0_avalon_master_readdata;                // mm_interconnect_0:framebuffer_sdram_0_avalon_master_readdata -> framebuffer_sdram_0:m0_readdata
	wire  [25:0] framebuffer_sdram_0_avalon_master_address;                 // framebuffer_sdram_0:m0_address -> mm_interconnect_0:framebuffer_sdram_0_avalon_master_address
	wire         framebuffer_sdram_0_avalon_master_read;                    // framebuffer_sdram_0:m0_read_n -> mm_interconnect_0:framebuffer_sdram_0_avalon_master_read
	wire   [1:0] framebuffer_sdram_0_avalon_master_byteenable;              // framebuffer_sdram_0:m0_byteenable_n -> mm_interconnect_0:framebuffer_sdram_0_avalon_master_byteenable
	wire         framebuffer_sdram_0_avalon_master_readdatavalid;           // mm_interconnect_0:framebuffer_sdram_0_avalon_master_readdatavalid -> framebuffer_sdram_0:m0_readdatavalid
	wire         framebuffer_sdram_0_avalon_master_write;                   // framebuffer_sdram_0:m0_write_n -> mm_interconnect_0:framebuffer_sdram_0_avalon_master_write
	wire  [15:0] framebuffer_sdram_0_avalon_master_writedata;               // framebuffer_sdram_0:m0_writedata -> mm_interconnect_0:framebuffer_sdram_0_avalon_master_writedata
	wire  [31:0] cpu_data_master_readdata;                                  // mm_interconnect_0:cpu_data_master_readdata -> cpu:d_readdata
	wire         cpu_data_master_waitrequest;                               // mm_interconnect_0:cpu_data_master_waitrequest -> cpu:d_waitrequest
	wire         cpu_data_master_debugaccess;                               // cpu:debug_mem_slave_debugaccess_to_roms -> mm_interconnect_0:cpu_data_master_debugaccess
	wire  [26:0] cpu_data_master_address;                                   // cpu:d_address -> mm_interconnect_0:cpu_data_master_address
	wire   [3:0] cpu_data_master_byteenable;                                // cpu:d_byteenable -> mm_interconnect_0:cpu_data_master_byteenable
	wire         cpu_data_master_read;                                      // cpu:d_read -> mm_interconnect_0:cpu_data_master_read
	wire         cpu_data_master_write;                                     // cpu:d_write -> mm_interconnect_0:cpu_data_master_write
	wire  [31:0] cpu_data_master_writedata;                                 // cpu:d_writedata -> mm_interconnect_0:cpu_data_master_writedata
	wire  [31:0] cpu_instruction_master_readdata;                           // mm_interconnect_0:cpu_instruction_master_readdata -> cpu:i_readdata
	wire         cpu_instruction_master_waitrequest;                        // mm_interconnect_0:cpu_instruction_master_waitrequest -> cpu:i_waitrequest
	wire  [26:0] cpu_instruction_master_address;                            // cpu:i_address -> mm_interconnect_0:cpu_instruction_master_address
	wire         cpu_instruction_master_read;                               // cpu:i_read -> mm_interconnect_0:cpu_instruction_master_read
	wire         mm_interconnect_0_new_sdram_controller_0_s1_chipselect;    // mm_interconnect_0:new_sdram_controller_0_s1_chipselect -> new_sdram_controller_0:az_cs
	wire  [15:0] mm_interconnect_0_new_sdram_controller_0_s1_readdata;      // new_sdram_controller_0:za_data -> mm_interconnect_0:new_sdram_controller_0_s1_readdata
	wire         mm_interconnect_0_new_sdram_controller_0_s1_waitrequest;   // new_sdram_controller_0:za_waitrequest -> mm_interconnect_0:new_sdram_controller_0_s1_waitrequest
	wire  [24:0] mm_interconnect_0_new_sdram_controller_0_s1_address;       // mm_interconnect_0:new_sdram_controller_0_s1_address -> new_sdram_controller_0:az_addr
	wire         mm_interconnect_0_new_sdram_controller_0_s1_read;          // mm_interconnect_0:new_sdram_controller_0_s1_read -> new_sdram_controller_0:az_rd_n
	wire   [1:0] mm_interconnect_0_new_sdram_controller_0_s1_byteenable;    // mm_interconnect_0:new_sdram_controller_0_s1_byteenable -> new_sdram_controller_0:az_be_n
	wire         mm_interconnect_0_new_sdram_controller_0_s1_readdatavalid; // new_sdram_controller_0:za_valid -> mm_interconnect_0:new_sdram_controller_0_s1_readdatavalid
	wire         mm_interconnect_0_new_sdram_controller_0_s1_write;         // mm_interconnect_0:new_sdram_controller_0_s1_write -> new_sdram_controller_0:az_wr_n
	wire  [15:0] mm_interconnect_0_new_sdram_controller_0_s1_writedata;     // mm_interconnect_0:new_sdram_controller_0_s1_writedata -> new_sdram_controller_0:az_data
	wire         mm_interconnect_0_jtag_uart_avalon_jtag_slave_chipselect;  // mm_interconnect_0:jtag_uart_avalon_jtag_slave_chipselect -> jtag_uart:av_chipselect
	wire  [31:0] mm_interconnect_0_jtag_uart_avalon_jtag_slave_readdata;    // jtag_uart:av_readdata -> mm_interconnect_0:jtag_uart_avalon_jtag_slave_readdata
	wire         mm_interconnect_0_jtag_uart_avalon_jtag_slave_waitrequest; // jtag_uart:av_waitrequest -> mm_interconnect_0:jtag_uart_avalon_jtag_slave_waitrequest
	wire   [0:0] mm_interconnect_0_jtag_uart_avalon_jtag_slave_address;     // mm_interconnect_0:jtag_uart_avalon_jtag_slave_address -> jtag_uart:av_address
	wire         mm_interconnect_0_jtag_uart_avalon_jtag_slave_read;        // mm_interconnect_0:jtag_uart_avalon_jtag_slave_read -> jtag_uart:av_read_n
	wire         mm_interconnect_0_jtag_uart_avalon_jtag_slave_write;       // mm_interconnect_0:jtag_uart_avalon_jtag_slave_write -> jtag_uart:av_write_n
	wire  [31:0] mm_interconnect_0_jtag_uart_avalon_jtag_slave_writedata;   // mm_interconnect_0:jtag_uart_avalon_jtag_slave_writedata -> jtag_uart:av_writedata
	wire  [31:0] mm_interconnect_0_cpu_debug_mem_slave_readdata;            // cpu:debug_mem_slave_readdata -> mm_interconnect_0:cpu_debug_mem_slave_readdata
	wire         mm_interconnect_0_cpu_debug_mem_slave_waitrequest;         // cpu:debug_mem_slave_waitrequest -> mm_interconnect_0:cpu_debug_mem_slave_waitrequest
	wire         mm_interconnect_0_cpu_debug_mem_slave_debugaccess;         // mm_interconnect_0:cpu_debug_mem_slave_debugaccess -> cpu:debug_mem_slave_debugaccess
	wire   [8:0] mm_interconnect_0_cpu_debug_mem_slave_address;             // mm_interconnect_0:cpu_debug_mem_slave_address -> cpu:debug_mem_slave_address
	wire         mm_interconnect_0_cpu_debug_mem_slave_read;                // mm_interconnect_0:cpu_debug_mem_slave_read -> cpu:debug_mem_slave_read
	wire   [3:0] mm_interconnect_0_cpu_debug_mem_slave_byteenable;          // mm_interconnect_0:cpu_debug_mem_slave_byteenable -> cpu:debug_mem_slave_byteenable
	wire         mm_interconnect_0_cpu_debug_mem_slave_write;               // mm_interconnect_0:cpu_debug_mem_slave_write -> cpu:debug_mem_slave_write
	wire  [31:0] mm_interconnect_0_cpu_debug_mem_slave_writedata;           // mm_interconnect_0:cpu_debug_mem_slave_writedata -> cpu:debug_mem_slave_writedata
	wire         mm_interconnect_0_i2c_avalon_0_i2c_chipselect;             // mm_interconnect_0:i2c_AVALON_0_i2c_chipselect -> i2c_AVALON_0:i2c_chipselect
	wire  [31:0] mm_interconnect_0_i2c_avalon_0_i2c_readdata;               // i2c_AVALON_0:i2c_readdata -> mm_interconnect_0:i2c_AVALON_0_i2c_readdata
	wire   [1:0] mm_interconnect_0_i2c_avalon_0_i2c_address;                // mm_interconnect_0:i2c_AVALON_0_i2c_address -> i2c_AVALON_0:i2c_address
	wire         mm_interconnect_0_i2c_avalon_0_i2c_write;                  // mm_interconnect_0:i2c_AVALON_0_i2c_write -> i2c_AVALON_0:i2c_write
	wire  [31:0] mm_interconnect_0_i2c_avalon_0_i2c_writedata;              // mm_interconnect_0:i2c_AVALON_0_i2c_writedata -> i2c_AVALON_0:i2c_writedata
	wire  [31:0] mm_interconnect_0_framebuffer_sdram_0_s0_readdata;         // framebuffer_sdram_0:s0_readdata -> mm_interconnect_0:framebuffer_sdram_0_s0_readdata
	wire   [0:0] mm_interconnect_0_framebuffer_sdram_0_s0_address;          // mm_interconnect_0:framebuffer_sdram_0_s0_address -> framebuffer_sdram_0:s0_address
	wire         mm_interconnect_0_framebuffer_sdram_0_s0_read;             // mm_interconnect_0:framebuffer_sdram_0_s0_read -> framebuffer_sdram_0:s0_read
	wire         mm_interconnect_0_framebuffer_sdram_0_s0_write;            // mm_interconnect_0:framebuffer_sdram_0_s0_write -> framebuffer_sdram_0:s0_write
	wire  [31:0] mm_interconnect_0_framebuffer_sdram_0_s0_writedata;        // mm_interconnect_0:framebuffer_sdram_0_s0_writedata -> framebuffer_sdram_0:s0_writedata
	wire         mm_interconnect_0_onchip_memory2_s1_chipselect;            // mm_interconnect_0:onchip_memory2_s1_chipselect -> onchip_memory2:chipselect
	wire  [31:0] mm_interconnect_0_onchip_memory2_s1_readdata;              // onchip_memory2:readdata -> mm_interconnect_0:onchip_memory2_s1_readdata
	wire  [15:0] mm_interconnect_0_onchip_memory2_s1_address;               // mm_interconnect_0:onchip_memory2_s1_address -> onchip_memory2:address
	wire   [3:0] mm_interconnect_0_onchip_memory2_s1_byteenable;            // mm_interconnect_0:onchip_memory2_s1_byteenable -> onchip_memory2:byteenable
	wire         mm_interconnect_0_onchip_memory2_s1_write;                 // mm_interconnect_0:onchip_memory2_s1_write -> onchip_memory2:write
	wire  [31:0] mm_interconnect_0_onchip_memory2_s1_writedata;             // mm_interconnect_0:onchip_memory2_s1_writedata -> onchip_memory2:writedata
	wire         mm_interconnect_0_onchip_memory2_s1_clken;                 // mm_interconnect_0:onchip_memory2_s1_clken -> onchip_memory2:clken
	wire         mm_interconnect_0_spi_avalon_sd_0_sd_chipselect;           // mm_interconnect_0:SPI_AVALON_SD_0_sd_chipselect -> SPI_AVALON_SD_0:sd_chipselect
	wire  [31:0] mm_interconnect_0_spi_avalon_sd_0_sd_readdata;             // SPI_AVALON_SD_0:sd_readdata -> mm_interconnect_0:SPI_AVALON_SD_0_sd_readdata
	wire   [1:0] mm_interconnect_0_spi_avalon_sd_0_sd_address;              // mm_interconnect_0:SPI_AVALON_SD_0_sd_address -> SPI_AVALON_SD_0:sd_address
	wire         mm_interconnect_0_spi_avalon_sd_0_sd_write;                // mm_interconnect_0:SPI_AVALON_SD_0_sd_write -> SPI_AVALON_SD_0:sd_write
	wire  [31:0] mm_interconnect_0_spi_avalon_sd_0_sd_writedata;            // mm_interconnect_0:SPI_AVALON_SD_0_sd_writedata -> SPI_AVALON_SD_0:sd_writedata
	wire         irq_mapper_receiver0_irq;                                  // jtag_uart:av_irq -> irq_mapper:receiver0_irq
	wire  [31:0] cpu_irq_irq;                                               // irq_mapper:sender_irq -> cpu:irq
	wire         rst_controller_reset_out_reset;                            // rst_controller:reset_out -> [SPI_AVALON_SD_0:reset, cpu:reset_n, framebuffer_sdram_0:rst, i2c_AVALON_0:reset, irq_mapper:reset, jtag_uart:rst_n, mm_interconnect_0:framebuffer_sdram_0_rst_reset_bridge_in_reset_reset, new_sdram_controller_0:reset_n, onchip_memory2:reset, rst_translator:in_reset]
	wire         rst_controller_reset_out_reset_req;                        // rst_controller:reset_req -> [cpu:reset_req, onchip_memory2:reset_req, rst_translator:reset_req_in]

	SPI_AVALON_SD spi_avalon_sd_0 (
		.clk           (pll_outclk0_clk),                                 //       clock.clk
		.reset         (rst_controller_reset_out_reset),                  //       reset.reset
		.sd_chipselect (mm_interconnect_0_spi_avalon_sd_0_sd_chipselect), //          sd.chipselect
		.sd_write      (mm_interconnect_0_spi_avalon_sd_0_sd_write),      //            .write
		.sd_address    (mm_interconnect_0_spi_avalon_sd_0_sd_address),    //            .address
		.sd_writedata  (mm_interconnect_0_spi_avalon_sd_0_sd_writedata),  //            .writedata
		.sd_readdata   (mm_interconnect_0_spi_avalon_sd_0_sd_readdata),   //            .readdata
		.sd_cs         (sd_sd_cs),                                        // conduit_end.sd_cs
		.sd_clk        (sd_sd_clk),                                       //            .sd_clk
		.sd_di         (sd_sd_di),                                        //            .sd_di
		.sd_do         (sd_sd_do)                                         //            .sd_do
	);

	DE1_SOC_NIOS_2_cpu cpu (
		.clk                                 (pll_outclk0_clk),                                   //                       clk.clk
		.reset_n                             (~rst_controller_reset_out_reset),                   //                     reset.reset_n
		.reset_req                           (rst_controller_reset_out_reset_req),                //                          .reset_req
		.d_address                           (cpu_data_master_address),                           //               data_master.address
		.d_byteenable                        (cpu_data_master_byteenable),                        //                          .byteenable
		.d_read                              (cpu_data_master_read),                              //                          .read
		.d_readdata                          (cpu_data_master_readdata),                          //                          .readdata
		.d_waitrequest                       (cpu_data_master_waitrequest),                       //                          .waitrequest
		.d_write                             (cpu_data_master_write),                             //                          .write
		.d_writedata                         (cpu_data_master_writedata),                         //                          .writedata
		.debug_mem_slave_debugaccess_to_roms (cpu_data_master_debugaccess),                       //                          .debugaccess
		.i_address                           (cpu_instruction_master_address),                    //        instruction_master.address
		.i_read                              (cpu_instruction_master_read),                       //                          .read
		.i_readdata                          (cpu_instruction_master_readdata),                   //                          .readdata
		.i_waitrequest                       (cpu_instruction_master_waitrequest),                //                          .waitrequest
		.irq                                 (cpu_irq_irq),                                       //                       irq.irq
		.debug_reset_request                 (),                                                  //       debug_reset_request.reset
		.debug_mem_slave_address             (mm_interconnect_0_cpu_debug_mem_slave_address),     //           debug_mem_slave.address
		.debug_mem_slave_byteenable          (mm_interconnect_0_cpu_debug_mem_slave_byteenable),  //                          .byteenable
		.debug_mem_slave_debugaccess         (mm_interconnect_0_cpu_debug_mem_slave_debugaccess), //                          .debugaccess
		.debug_mem_slave_read                (mm_interconnect_0_cpu_debug_mem_slave_read),        //                          .read
		.debug_mem_slave_readdata            (mm_interconnect_0_cpu_debug_mem_slave_readdata),    //                          .readdata
		.debug_mem_slave_waitrequest         (mm_interconnect_0_cpu_debug_mem_slave_waitrequest), //                          .waitrequest
		.debug_mem_slave_write               (mm_interconnect_0_cpu_debug_mem_slave_write),       //                          .write
		.debug_mem_slave_writedata           (mm_interconnect_0_cpu_debug_mem_slave_writedata),   //                          .writedata
		.dummy_ci_port                       ()                                                   // custom_instruction_master.readra
	);

	framebuffer_arbiter framebuffer_sdram_0 (
		.clk                 (pll_outclk0_clk),                                    //         clock.clk
		.s0_address          (mm_interconnect_0_framebuffer_sdram_0_s0_address),   //            s0.address
		.s0_read             (mm_interconnect_0_framebuffer_sdram_0_s0_read),      //              .read
		.s0_write            (mm_interconnect_0_framebuffer_sdram_0_s0_write),     //              .write
		.s0_writedata        (mm_interconnect_0_framebuffer_sdram_0_s0_writedata), //              .writedata
		.s0_readdata         (mm_interconnect_0_framebuffer_sdram_0_s0_readdata),  //              .readdata
		.m0_waitrequest      (framebuffer_sdram_0_avalon_master_waitrequest),      // avalon_master.waitrequest
		.m0_readdatavalid    (framebuffer_sdram_0_avalon_master_readdatavalid),    //              .readdatavalid
		.m0_readdata         (framebuffer_sdram_0_avalon_master_readdata),         //              .readdata
		.m0_address          (framebuffer_sdram_0_avalon_master_address),          //              .address
		.m0_read_n           (framebuffer_sdram_0_avalon_master_read),             //              .read_n
		.m0_chipselect       (framebuffer_sdram_0_avalon_master_chipselect),       //              .chipselect
		.m0_byteenable_n     (framebuffer_sdram_0_avalon_master_byteenable),       //              .byteenable_n
		.m0_write_n          (framebuffer_sdram_0_avalon_master_write),            //              .write_n
		.m0_writedata        (framebuffer_sdram_0_avalon_master_writedata),        //              .writedata
		.rst                 (rst_controller_reset_out_reset),                     //           rst.reset
		.export_read_clk     (pixel_read_clk),                                     //        export.read_clk
		.export_as0_ready    (pixel_ready),                                        //              .ready
		.export_as0_valid    (pixel_valid),                                        //              .valid
		.export_as0_readdata (pixel_readdata),                                     //              .readdata
		.export_frame_sync   (pixel_frame_sync)                                    //              .frame_sync
	);

	I2C_AVALON i2c_avalon_0 (
		.clk            (pll_outclk0_clk),                               //       clock.clk
		.reset          (rst_controller_reset_out_reset),                //       reset.reset
		.i2c_chipselect (mm_interconnect_0_i2c_avalon_0_i2c_chipselect), //         i2c.chipselect
		.i2c_write      (mm_interconnect_0_i2c_avalon_0_i2c_write),      //            .write
		.i2c_address    (mm_interconnect_0_i2c_avalon_0_i2c_address),    //            .address
		.i2c_writedata  (mm_interconnect_0_i2c_avalon_0_i2c_writedata),  //            .writedata
		.i2c_readdata   (mm_interconnect_0_i2c_avalon_0_i2c_readdata),   //            .readdata
		.i2c_reset      (i2c_rst),                                       // conduit_end.rst
		.i2c_sda        (i2c_sda),                                       //            .sda
		.i2c_sclk       (i2c_sclk)                                       //            .sclk
	);

	DE1_SOC_NIOS_2_jtag_uart jtag_uart (
		.clk            (pll_outclk0_clk),                                           //               clk.clk
		.rst_n          (~rst_controller_reset_out_reset),                           //             reset.reset_n
		.av_chipselect  (mm_interconnect_0_jtag_uart_avalon_jtag_slave_chipselect),  // avalon_jtag_slave.chipselect
		.av_address     (mm_interconnect_0_jtag_uart_avalon_jtag_slave_address),     //                  .address
		.av_read_n      (~mm_interconnect_0_jtag_uart_avalon_jtag_slave_read),       //                  .read_n
		.av_readdata    (mm_interconnect_0_jtag_uart_avalon_jtag_slave_readdata),    //                  .readdata
		.av_write_n     (~mm_interconnect_0_jtag_uart_avalon_jtag_slave_write),      //                  .write_n
		.av_writedata   (mm_interconnect_0_jtag_uart_avalon_jtag_slave_writedata),   //                  .writedata
		.av_waitrequest (mm_interconnect_0_jtag_uart_avalon_jtag_slave_waitrequest), //                  .waitrequest
		.av_irq         (irq_mapper_receiver0_irq)                                   //               irq.irq
	);

	DE1_SOC_NIOS_2_new_sdram_controller_0 new_sdram_controller_0 (
		.clk            (pll_outclk0_clk),                                           //   clk.clk
		.reset_n        (~rst_controller_reset_out_reset),                           // reset.reset_n
		.az_addr        (mm_interconnect_0_new_sdram_controller_0_s1_address),       //    s1.address
		.az_be_n        (~mm_interconnect_0_new_sdram_controller_0_s1_byteenable),   //      .byteenable_n
		.az_cs          (mm_interconnect_0_new_sdram_controller_0_s1_chipselect),    //      .chipselect
		.az_data        (mm_interconnect_0_new_sdram_controller_0_s1_writedata),     //      .writedata
		.az_rd_n        (~mm_interconnect_0_new_sdram_controller_0_s1_read),         //      .read_n
		.az_wr_n        (~mm_interconnect_0_new_sdram_controller_0_s1_write),        //      .write_n
		.za_data        (mm_interconnect_0_new_sdram_controller_0_s1_readdata),      //      .readdata
		.za_valid       (mm_interconnect_0_new_sdram_controller_0_s1_readdatavalid), //      .readdatavalid
		.za_waitrequest (mm_interconnect_0_new_sdram_controller_0_s1_waitrequest),   //      .waitrequest
		.zs_addr        (new_sdram_controller_0_wire_addr),                          //  wire.export
		.zs_ba          (new_sdram_controller_0_wire_ba),                            //      .export
		.zs_cas_n       (new_sdram_controller_0_wire_cas_n),                         //      .export
		.zs_cke         (new_sdram_controller_0_wire_cke),                           //      .export
		.zs_cs_n        (new_sdram_controller_0_wire_cs_n),                          //      .export
		.zs_dq          (new_sdram_controller_0_wire_dq),                            //      .export
		.zs_dqm         (new_sdram_controller_0_wire_dqm),                           //      .export
		.zs_ras_n       (new_sdram_controller_0_wire_ras_n),                         //      .export
		.zs_we_n        (new_sdram_controller_0_wire_we_n)                           //      .export
	);

	DE1_SOC_NIOS_2_onchip_memory2 onchip_memory2 (
		.clk        (pll_outclk0_clk),                                //   clk1.clk
		.address    (mm_interconnect_0_onchip_memory2_s1_address),    //     s1.address
		.clken      (mm_interconnect_0_onchip_memory2_s1_clken),      //       .clken
		.chipselect (mm_interconnect_0_onchip_memory2_s1_chipselect), //       .chipselect
		.write      (mm_interconnect_0_onchip_memory2_s1_write),      //       .write
		.readdata   (mm_interconnect_0_onchip_memory2_s1_readdata),   //       .readdata
		.writedata  (mm_interconnect_0_onchip_memory2_s1_writedata),  //       .writedata
		.byteenable (mm_interconnect_0_onchip_memory2_s1_byteenable), //       .byteenable
		.reset      (rst_controller_reset_out_reset),                 // reset1.reset
		.reset_req  (rst_controller_reset_out_reset_req)              //       .reset_req
	);

	DE1_SOC_NIOS_2_pll pll (
		.refclk   (clk_clk),         //  refclk.clk
		.rst      (~reset_reset_n),  //   reset.reset
		.outclk_0 (pll_outclk0_clk), // outclk0.clk
		.outclk_1 (sdram_clk_clk),   // outclk1.clk
		.locked   ()                 // (terminated)
	);

	DE1_SOC_NIOS_2_pll_I2C pll_i2c (
		.refclk   (clk_clk),         //  refclk.clk
		.rst      (~reset_reset_n),  //   reset.reset
		.outclk_0 (clock_6400k_clk), // outclk0.clk
		.outclk_1 (clock_23m_clk),   // outclk1.clk
		.locked   ()                 // (terminated)
	);

	DE1_SOC_NIOS_2_mm_interconnect_0 mm_interconnect_0 (
		.pll_outclk0_clk                                     (pll_outclk0_clk),                                           //                                   pll_outclk0.clk
		.framebuffer_sdram_0_rst_reset_bridge_in_reset_reset (rst_controller_reset_out_reset),                            // framebuffer_sdram_0_rst_reset_bridge_in_reset.reset
		.cpu_data_master_address                             (cpu_data_master_address),                                   //                               cpu_data_master.address
		.cpu_data_master_waitrequest                         (cpu_data_master_waitrequest),                               //                                              .waitrequest
		.cpu_data_master_byteenable                          (cpu_data_master_byteenable),                                //                                              .byteenable
		.cpu_data_master_read                                (cpu_data_master_read),                                      //                                              .read
		.cpu_data_master_readdata                            (cpu_data_master_readdata),                                  //                                              .readdata
		.cpu_data_master_write                               (cpu_data_master_write),                                     //                                              .write
		.cpu_data_master_writedata                           (cpu_data_master_writedata),                                 //                                              .writedata
		.cpu_data_master_debugaccess                         (cpu_data_master_debugaccess),                               //                                              .debugaccess
		.cpu_instruction_master_address                      (cpu_instruction_master_address),                            //                        cpu_instruction_master.address
		.cpu_instruction_master_waitrequest                  (cpu_instruction_master_waitrequest),                        //                                              .waitrequest
		.cpu_instruction_master_read                         (cpu_instruction_master_read),                               //                                              .read
		.cpu_instruction_master_readdata                     (cpu_instruction_master_readdata),                           //                                              .readdata
		.framebuffer_sdram_0_avalon_master_address           (framebuffer_sdram_0_avalon_master_address),                 //             framebuffer_sdram_0_avalon_master.address
		.framebuffer_sdram_0_avalon_master_waitrequest       (framebuffer_sdram_0_avalon_master_waitrequest),             //                                              .waitrequest
		.framebuffer_sdram_0_avalon_master_byteenable        (~framebuffer_sdram_0_avalon_master_byteenable),             //                                              .byteenable
		.framebuffer_sdram_0_avalon_master_chipselect        (framebuffer_sdram_0_avalon_master_chipselect),              //                                              .chipselect
		.framebuffer_sdram_0_avalon_master_read              (~framebuffer_sdram_0_avalon_master_read),                   //                                              .read
		.framebuffer_sdram_0_avalon_master_readdata          (framebuffer_sdram_0_avalon_master_readdata),                //                                              .readdata
		.framebuffer_sdram_0_avalon_master_readdatavalid     (framebuffer_sdram_0_avalon_master_readdatavalid),           //                                              .readdatavalid
		.framebuffer_sdram_0_avalon_master_write             (~framebuffer_sdram_0_avalon_master_write),                  //                                              .write
		.framebuffer_sdram_0_avalon_master_writedata         (framebuffer_sdram_0_avalon_master_writedata),               //                                              .writedata
		.cpu_debug_mem_slave_address                         (mm_interconnect_0_cpu_debug_mem_slave_address),             //                           cpu_debug_mem_slave.address
		.cpu_debug_mem_slave_write                           (mm_interconnect_0_cpu_debug_mem_slave_write),               //                                              .write
		.cpu_debug_mem_slave_read                            (mm_interconnect_0_cpu_debug_mem_slave_read),                //                                              .read
		.cpu_debug_mem_slave_readdata                        (mm_interconnect_0_cpu_debug_mem_slave_readdata),            //                                              .readdata
		.cpu_debug_mem_slave_writedata                       (mm_interconnect_0_cpu_debug_mem_slave_writedata),           //                                              .writedata
		.cpu_debug_mem_slave_byteenable                      (mm_interconnect_0_cpu_debug_mem_slave_byteenable),          //                                              .byteenable
		.cpu_debug_mem_slave_waitrequest                     (mm_interconnect_0_cpu_debug_mem_slave_waitrequest),         //                                              .waitrequest
		.cpu_debug_mem_slave_debugaccess                     (mm_interconnect_0_cpu_debug_mem_slave_debugaccess),         //                                              .debugaccess
		.framebuffer_sdram_0_s0_address                      (mm_interconnect_0_framebuffer_sdram_0_s0_address),          //                        framebuffer_sdram_0_s0.address
		.framebuffer_sdram_0_s0_write                        (mm_interconnect_0_framebuffer_sdram_0_s0_write),            //                                              .write
		.framebuffer_sdram_0_s0_read                         (mm_interconnect_0_framebuffer_sdram_0_s0_read),             //                                              .read
		.framebuffer_sdram_0_s0_readdata                     (mm_interconnect_0_framebuffer_sdram_0_s0_readdata),         //                                              .readdata
		.framebuffer_sdram_0_s0_writedata                    (mm_interconnect_0_framebuffer_sdram_0_s0_writedata),        //                                              .writedata
		.i2c_AVALON_0_i2c_address                            (mm_interconnect_0_i2c_avalon_0_i2c_address),                //                              i2c_AVALON_0_i2c.address
		.i2c_AVALON_0_i2c_write                              (mm_interconnect_0_i2c_avalon_0_i2c_write),                  //                                              .write
		.i2c_AVALON_0_i2c_readdata                           (mm_interconnect_0_i2c_avalon_0_i2c_readdata),               //                                              .readdata
		.i2c_AVALON_0_i2c_writedata                          (mm_interconnect_0_i2c_avalon_0_i2c_writedata),              //                                              .writedata
		.i2c_AVALON_0_i2c_chipselect                         (mm_interconnect_0_i2c_avalon_0_i2c_chipselect),             //                                              .chipselect
		.jtag_uart_avalon_jtag_slave_address                 (mm_interconnect_0_jtag_uart_avalon_jtag_slave_address),     //                   jtag_uart_avalon_jtag_slave.address
		.jtag_uart_avalon_jtag_slave_write                   (mm_interconnect_0_jtag_uart_avalon_jtag_slave_write),       //                                              .write
		.jtag_uart_avalon_jtag_slave_read                    (mm_interconnect_0_jtag_uart_avalon_jtag_slave_read),        //                                              .read
		.jtag_uart_avalon_jtag_slave_readdata                (mm_interconnect_0_jtag_uart_avalon_jtag_slave_readdata),    //                                              .readdata
		.jtag_uart_avalon_jtag_slave_writedata               (mm_interconnect_0_jtag_uart_avalon_jtag_slave_writedata),   //                                              .writedata
		.jtag_uart_avalon_jtag_slave_waitrequest             (mm_interconnect_0_jtag_uart_avalon_jtag_slave_waitrequest), //                                              .waitrequest
		.jtag_uart_avalon_jtag_slave_chipselect              (mm_interconnect_0_jtag_uart_avalon_jtag_slave_chipselect),  //                                              .chipselect
		.new_sdram_controller_0_s1_address                   (mm_interconnect_0_new_sdram_controller_0_s1_address),       //                     new_sdram_controller_0_s1.address
		.new_sdram_controller_0_s1_write                     (mm_interconnect_0_new_sdram_controller_0_s1_write),         //                                              .write
		.new_sdram_controller_0_s1_read                      (mm_interconnect_0_new_sdram_controller_0_s1_read),          //                                              .read
		.new_sdram_controller_0_s1_readdata                  (mm_interconnect_0_new_sdram_controller_0_s1_readdata),      //                                              .readdata
		.new_sdram_controller_0_s1_writedata                 (mm_interconnect_0_new_sdram_controller_0_s1_writedata),     //                                              .writedata
		.new_sdram_controller_0_s1_byteenable                (mm_interconnect_0_new_sdram_controller_0_s1_byteenable),    //                                              .byteenable
		.new_sdram_controller_0_s1_readdatavalid             (mm_interconnect_0_new_sdram_controller_0_s1_readdatavalid), //                                              .readdatavalid
		.new_sdram_controller_0_s1_waitrequest               (mm_interconnect_0_new_sdram_controller_0_s1_waitrequest),   //                                              .waitrequest
		.new_sdram_controller_0_s1_chipselect                (mm_interconnect_0_new_sdram_controller_0_s1_chipselect),    //                                              .chipselect
		.onchip_memory2_s1_address                           (mm_interconnect_0_onchip_memory2_s1_address),               //                             onchip_memory2_s1.address
		.onchip_memory2_s1_write                             (mm_interconnect_0_onchip_memory2_s1_write),                 //                                              .write
		.onchip_memory2_s1_readdata                          (mm_interconnect_0_onchip_memory2_s1_readdata),              //                                              .readdata
		.onchip_memory2_s1_writedata                         (mm_interconnect_0_onchip_memory2_s1_writedata),             //                                              .writedata
		.onchip_memory2_s1_byteenable                        (mm_interconnect_0_onchip_memory2_s1_byteenable),            //                                              .byteenable
		.onchip_memory2_s1_chipselect                        (mm_interconnect_0_onchip_memory2_s1_chipselect),            //                                              .chipselect
		.onchip_memory2_s1_clken                             (mm_interconnect_0_onchip_memory2_s1_clken),                 //                                              .clken
		.SPI_AVALON_SD_0_sd_address                          (mm_interconnect_0_spi_avalon_sd_0_sd_address),              //                            SPI_AVALON_SD_0_sd.address
		.SPI_AVALON_SD_0_sd_write                            (mm_interconnect_0_spi_avalon_sd_0_sd_write),                //                                              .write
		.SPI_AVALON_SD_0_sd_readdata                         (mm_interconnect_0_spi_avalon_sd_0_sd_readdata),             //                                              .readdata
		.SPI_AVALON_SD_0_sd_writedata                        (mm_interconnect_0_spi_avalon_sd_0_sd_writedata),            //                                              .writedata
		.SPI_AVALON_SD_0_sd_chipselect                       (mm_interconnect_0_spi_avalon_sd_0_sd_chipselect)            //                                              .chipselect
	);

	DE1_SOC_NIOS_2_irq_mapper irq_mapper (
		.clk           (pll_outclk0_clk),                //       clk.clk
		.reset         (rst_controller_reset_out_reset), // clk_reset.reset
		.receiver0_irq (irq_mapper_receiver0_irq),       // receiver0.irq
		.sender_irq    (cpu_irq_irq)                     //    sender.irq
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (1),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller (
		.reset_in0      (~reset_reset_n),                     // reset_in0.reset
		.clk            (pll_outclk0_clk),                    //       clk.clk
		.reset_out      (rst_controller_reset_out_reset),     // reset_out.reset
		.reset_req      (rst_controller_reset_out_reset_req), //          .reset_req
		.reset_req_in0  (1'b0),                               // (terminated)
		.reset_in1      (1'b0),                               // (terminated)
		.reset_req_in1  (1'b0),                               // (terminated)
		.reset_in2      (1'b0),                               // (terminated)
		.reset_req_in2  (1'b0),                               // (terminated)
		.reset_in3      (1'b0),                               // (terminated)
		.reset_req_in3  (1'b0),                               // (terminated)
		.reset_in4      (1'b0),                               // (terminated)
		.reset_req_in4  (1'b0),                               // (terminated)
		.reset_in5      (1'b0),                               // (terminated)
		.reset_req_in5  (1'b0),                               // (terminated)
		.reset_in6      (1'b0),                               // (terminated)
		.reset_req_in6  (1'b0),                               // (terminated)
		.reset_in7      (1'b0),                               // (terminated)
		.reset_req_in7  (1'b0),                               // (terminated)
		.reset_in8      (1'b0),                               // (terminated)
		.reset_req_in8  (1'b0),                               // (terminated)
		.reset_in9      (1'b0),                               // (terminated)
		.reset_req_in9  (1'b0),                               // (terminated)
		.reset_in10     (1'b0),                               // (terminated)
		.reset_req_in10 (1'b0),                               // (terminated)
		.reset_in11     (1'b0),                               // (terminated)
		.reset_req_in11 (1'b0),                               // (terminated)
		.reset_in12     (1'b0),                               // (terminated)
		.reset_req_in12 (1'b0),                               // (terminated)
		.reset_in13     (1'b0),                               // (terminated)
		.reset_req_in13 (1'b0),                               // (terminated)
		.reset_in14     (1'b0),                               // (terminated)
		.reset_req_in14 (1'b0),                               // (terminated)
		.reset_in15     (1'b0),                               // (terminated)
		.reset_req_in15 (1'b0)                                // (terminated)
	);

endmodule
