// DE1_SOC_NIOS_2.v

// Generated using ACDS version 15.0 145

`timescale 1 ps / 1 ps
module DE1_SOC_NIOS_2 (
		input  wire        clk_clk,                           //                         clk.clk
		output wire        i2c_rst,                           //                         i2c.rst
		inout  wire        i2c_sda,                           //                            .sda
		inout  wire        i2c_sclk,                          //                            .sclk
		output wire        lcd_lcd_cs,                        //                         lcd.lcd_cs
		output wire [23:0] lcd_lcd_data,                      //                            .lcd_data
		output wire        lcd_lcd_dc,                        //                            .lcd_dc
		output wire        lcd_lcd_rst,                       //                            .lcd_rst
		output wire        lcd_lcd_wr,                        //                            .lcd_wr
		output wire [12:0] new_sdram_controller_0_wire_addr,  // new_sdram_controller_0_wire.addr
		output wire [1:0]  new_sdram_controller_0_wire_ba,    //                            .ba
		output wire        new_sdram_controller_0_wire_cas_n, //                            .cas_n
		output wire        new_sdram_controller_0_wire_cke,   //                            .cke
		output wire        new_sdram_controller_0_wire_cs_n,  //                            .cs_n
		inout  wire [15:0] new_sdram_controller_0_wire_dq,    //                            .dq
		output wire [1:0]  new_sdram_controller_0_wire_dqm,   //                            .dqm
		output wire        new_sdram_controller_0_wire_ras_n, //                            .ras_n
		output wire        new_sdram_controller_0_wire_we_n,  //                            .we_n
		input  wire        reset_reset_n,                     //                       reset.reset_n
		output wire        sd_sd_cs,                          //                          sd.sd_cs
		output wire        sd_sd_clk,                         //                            .sd_clk
		output wire        sd_sd_di,                          //                            .sd_di
		input  wire        sd_sd_do,                          //                            .sd_do
		output wire        sdram_clk_clk                      //                   sdram_clk.clk
	);

	wire         pll_outclk0_clk;                                           // pll:outclk_0 -> [SPI_AVALON_SD_0:clk, cpu:clk, i2c_AVALON_0:clk, irq_mapper:clk, irq_synchronizer:sender_clk, irq_synchronizer_001:sender_clk, jtag_uart:clk, mm_interconnect_0:pll_outclk0_clk, new_sdram_controller_0:clk, onchip_memory2:clk, rst_controller_001:clk]
	wire         lcdframebuffer_0_avalon_master_chipselect;                 // LCDFrameBuffer_0:m0_chipselect -> mm_interconnect_0:LCDFrameBuffer_0_avalon_master_chipselect
	wire         lcdframebuffer_0_avalon_master_waitrequest;                // mm_interconnect_0:LCDFrameBuffer_0_avalon_master_waitrequest -> LCDFrameBuffer_0:m0_waitrequest
	wire  [15:0] lcdframebuffer_0_avalon_master_readdata;                   // mm_interconnect_0:LCDFrameBuffer_0_avalon_master_readdata -> LCDFrameBuffer_0:m0_readdata
	wire  [25:0] lcdframebuffer_0_avalon_master_address;                    // LCDFrameBuffer_0:m0_address -> mm_interconnect_0:LCDFrameBuffer_0_avalon_master_address
	wire   [1:0] lcdframebuffer_0_avalon_master_byteenable;                 // LCDFrameBuffer_0:m0_byteenable_n -> mm_interconnect_0:LCDFrameBuffer_0_avalon_master_byteenable
	wire         lcdframebuffer_0_avalon_master_read;                       // LCDFrameBuffer_0:m0_read_n -> mm_interconnect_0:LCDFrameBuffer_0_avalon_master_read
	wire         lcdframebuffer_0_avalon_master_readdatavalid;              // mm_interconnect_0:LCDFrameBuffer_0_avalon_master_readdatavalid -> LCDFrameBuffer_0:m0_readdatavalid
	wire  [15:0] lcdframebuffer_0_avalon_master_writedata;                  // LCDFrameBuffer_0:m0_writedata -> mm_interconnect_0:LCDFrameBuffer_0_avalon_master_writedata
	wire         lcdframebuffer_0_avalon_master_write;                      // LCDFrameBuffer_0:m0_write_n -> mm_interconnect_0:LCDFrameBuffer_0_avalon_master_write
	wire  [31:0] cpu_data_master_readdata;                                  // mm_interconnect_0:cpu_data_master_readdata -> cpu:d_readdata
	wire         cpu_data_master_waitrequest;                               // mm_interconnect_0:cpu_data_master_waitrequest -> cpu:d_waitrequest
	wire         cpu_data_master_debugaccess;                               // cpu:debug_mem_slave_debugaccess_to_roms -> mm_interconnect_0:cpu_data_master_debugaccess
	wire  [26:0] cpu_data_master_address;                                   // cpu:d_address -> mm_interconnect_0:cpu_data_master_address
	wire   [3:0] cpu_data_master_byteenable;                                // cpu:d_byteenable -> mm_interconnect_0:cpu_data_master_byteenable
	wire         cpu_data_master_read;                                      // cpu:d_read -> mm_interconnect_0:cpu_data_master_read
	wire         cpu_data_master_write;                                     // cpu:d_write -> mm_interconnect_0:cpu_data_master_write
	wire  [31:0] cpu_data_master_writedata;                                 // cpu:d_writedata -> mm_interconnect_0:cpu_data_master_writedata
	wire         dma_0_read_master_chipselect;                              // dma_0:read_chipselect -> mm_interconnect_0:dma_0_read_master_chipselect
	wire  [15:0] dma_0_read_master_readdata;                                // mm_interconnect_0:dma_0_read_master_readdata -> dma_0:read_readdata
	wire         dma_0_read_master_waitrequest;                             // mm_interconnect_0:dma_0_read_master_waitrequest -> dma_0:read_waitrequest
	wire  [25:0] dma_0_read_master_address;                                 // dma_0:read_address -> mm_interconnect_0:dma_0_read_master_address
	wire         dma_0_read_master_read;                                    // dma_0:read_read_n -> mm_interconnect_0:dma_0_read_master_read
	wire         dma_0_read_master_readdatavalid;                           // mm_interconnect_0:dma_0_read_master_readdatavalid -> dma_0:read_readdatavalid
	wire         dma_0_write_master_chipselect;                             // dma_0:write_chipselect -> mm_interconnect_0:dma_0_write_master_chipselect
	wire         dma_0_write_master_waitrequest;                            // mm_interconnect_0:dma_0_write_master_waitrequest -> dma_0:write_waitrequest
	wire  [25:0] dma_0_write_master_address;                                // dma_0:write_address -> mm_interconnect_0:dma_0_write_master_address
	wire   [1:0] dma_0_write_master_byteenable;                             // dma_0:write_byteenable -> mm_interconnect_0:dma_0_write_master_byteenable
	wire         dma_0_write_master_write;                                  // dma_0:write_write_n -> mm_interconnect_0:dma_0_write_master_write
	wire  [15:0] dma_0_write_master_writedata;                              // dma_0:write_writedata -> mm_interconnect_0:dma_0_write_master_writedata
	wire  [31:0] cpu_instruction_master_readdata;                           // mm_interconnect_0:cpu_instruction_master_readdata -> cpu:i_readdata
	wire         cpu_instruction_master_waitrequest;                        // mm_interconnect_0:cpu_instruction_master_waitrequest -> cpu:i_waitrequest
	wire  [26:0] cpu_instruction_master_address;                            // cpu:i_address -> mm_interconnect_0:cpu_instruction_master_address
	wire         cpu_instruction_master_read;                               // cpu:i_read -> mm_interconnect_0:cpu_instruction_master_read
	wire         mm_interconnect_0_new_sdram_controller_0_s1_chipselect;    // mm_interconnect_0:new_sdram_controller_0_s1_chipselect -> new_sdram_controller_0:az_cs
	wire  [15:0] mm_interconnect_0_new_sdram_controller_0_s1_readdata;      // new_sdram_controller_0:za_data -> mm_interconnect_0:new_sdram_controller_0_s1_readdata
	wire         mm_interconnect_0_new_sdram_controller_0_s1_waitrequest;   // new_sdram_controller_0:za_waitrequest -> mm_interconnect_0:new_sdram_controller_0_s1_waitrequest
	wire  [24:0] mm_interconnect_0_new_sdram_controller_0_s1_address;       // mm_interconnect_0:new_sdram_controller_0_s1_address -> new_sdram_controller_0:az_addr
	wire         mm_interconnect_0_new_sdram_controller_0_s1_read;          // mm_interconnect_0:new_sdram_controller_0_s1_read -> new_sdram_controller_0:az_rd_n
	wire   [1:0] mm_interconnect_0_new_sdram_controller_0_s1_byteenable;    // mm_interconnect_0:new_sdram_controller_0_s1_byteenable -> new_sdram_controller_0:az_be_n
	wire         mm_interconnect_0_new_sdram_controller_0_s1_readdatavalid; // new_sdram_controller_0:za_valid -> mm_interconnect_0:new_sdram_controller_0_s1_readdatavalid
	wire         mm_interconnect_0_new_sdram_controller_0_s1_write;         // mm_interconnect_0:new_sdram_controller_0_s1_write -> new_sdram_controller_0:az_wr_n
	wire  [15:0] mm_interconnect_0_new_sdram_controller_0_s1_writedata;     // mm_interconnect_0:new_sdram_controller_0_s1_writedata -> new_sdram_controller_0:az_data
	wire         mm_interconnect_0_jtag_uart_avalon_jtag_slave_chipselect;  // mm_interconnect_0:jtag_uart_avalon_jtag_slave_chipselect -> jtag_uart:av_chipselect
	wire  [31:0] mm_interconnect_0_jtag_uart_avalon_jtag_slave_readdata;    // jtag_uart:av_readdata -> mm_interconnect_0:jtag_uart_avalon_jtag_slave_readdata
	wire         mm_interconnect_0_jtag_uart_avalon_jtag_slave_waitrequest; // jtag_uart:av_waitrequest -> mm_interconnect_0:jtag_uart_avalon_jtag_slave_waitrequest
	wire   [0:0] mm_interconnect_0_jtag_uart_avalon_jtag_slave_address;     // mm_interconnect_0:jtag_uart_avalon_jtag_slave_address -> jtag_uart:av_address
	wire         mm_interconnect_0_jtag_uart_avalon_jtag_slave_read;        // mm_interconnect_0:jtag_uart_avalon_jtag_slave_read -> jtag_uart:av_read_n
	wire         mm_interconnect_0_jtag_uart_avalon_jtag_slave_write;       // mm_interconnect_0:jtag_uart_avalon_jtag_slave_write -> jtag_uart:av_write_n
	wire  [31:0] mm_interconnect_0_jtag_uart_avalon_jtag_slave_writedata;   // mm_interconnect_0:jtag_uart_avalon_jtag_slave_writedata -> jtag_uart:av_writedata
	wire         mm_interconnect_0_dma_0_control_port_slave_chipselect;     // mm_interconnect_0:dma_0_control_port_slave_chipselect -> dma_0:dma_ctl_chipselect
	wire  [25:0] mm_interconnect_0_dma_0_control_port_slave_readdata;       // dma_0:dma_ctl_readdata -> mm_interconnect_0:dma_0_control_port_slave_readdata
	wire   [2:0] mm_interconnect_0_dma_0_control_port_slave_address;        // mm_interconnect_0:dma_0_control_port_slave_address -> dma_0:dma_ctl_address
	wire         mm_interconnect_0_dma_0_control_port_slave_write;          // mm_interconnect_0:dma_0_control_port_slave_write -> dma_0:dma_ctl_write_n
	wire  [25:0] mm_interconnect_0_dma_0_control_port_slave_writedata;      // mm_interconnect_0:dma_0_control_port_slave_writedata -> dma_0:dma_ctl_writedata
	wire  [31:0] mm_interconnect_0_cpu_debug_mem_slave_readdata;            // cpu:debug_mem_slave_readdata -> mm_interconnect_0:cpu_debug_mem_slave_readdata
	wire         mm_interconnect_0_cpu_debug_mem_slave_waitrequest;         // cpu:debug_mem_slave_waitrequest -> mm_interconnect_0:cpu_debug_mem_slave_waitrequest
	wire         mm_interconnect_0_cpu_debug_mem_slave_debugaccess;         // mm_interconnect_0:cpu_debug_mem_slave_debugaccess -> cpu:debug_mem_slave_debugaccess
	wire   [8:0] mm_interconnect_0_cpu_debug_mem_slave_address;             // mm_interconnect_0:cpu_debug_mem_slave_address -> cpu:debug_mem_slave_address
	wire         mm_interconnect_0_cpu_debug_mem_slave_read;                // mm_interconnect_0:cpu_debug_mem_slave_read -> cpu:debug_mem_slave_read
	wire   [3:0] mm_interconnect_0_cpu_debug_mem_slave_byteenable;          // mm_interconnect_0:cpu_debug_mem_slave_byteenable -> cpu:debug_mem_slave_byteenable
	wire         mm_interconnect_0_cpu_debug_mem_slave_write;               // mm_interconnect_0:cpu_debug_mem_slave_write -> cpu:debug_mem_slave_write
	wire  [31:0] mm_interconnect_0_cpu_debug_mem_slave_writedata;           // mm_interconnect_0:cpu_debug_mem_slave_writedata -> cpu:debug_mem_slave_writedata
	wire         mm_interconnect_0_i2c_avalon_0_i2c_chipselect;             // mm_interconnect_0:i2c_AVALON_0_i2c_chipselect -> i2c_AVALON_0:i2c_chipselect
	wire  [31:0] mm_interconnect_0_i2c_avalon_0_i2c_readdata;               // i2c_AVALON_0:i2c_readdata -> mm_interconnect_0:i2c_AVALON_0_i2c_readdata
	wire   [1:0] mm_interconnect_0_i2c_avalon_0_i2c_address;                // mm_interconnect_0:i2c_AVALON_0_i2c_address -> i2c_AVALON_0:i2c_address
	wire         mm_interconnect_0_i2c_avalon_0_i2c_write;                  // mm_interconnect_0:i2c_AVALON_0_i2c_write -> i2c_AVALON_0:i2c_write
	wire  [31:0] mm_interconnect_0_i2c_avalon_0_i2c_writedata;              // mm_interconnect_0:i2c_AVALON_0_i2c_writedata -> i2c_AVALON_0:i2c_writedata
	wire         mm_interconnect_0_lcdframebuffer_0_s0_chipselect;          // mm_interconnect_0:LCDFrameBuffer_0_s0_chipselect -> LCDFrameBuffer_0:s0_chipselect
	wire  [31:0] mm_interconnect_0_lcdframebuffer_0_s0_readdata;            // LCDFrameBuffer_0:s0_readdata -> mm_interconnect_0:LCDFrameBuffer_0_s0_readdata
	wire   [1:0] mm_interconnect_0_lcdframebuffer_0_s0_address;             // mm_interconnect_0:LCDFrameBuffer_0_s0_address -> LCDFrameBuffer_0:s0_address
	wire         mm_interconnect_0_lcdframebuffer_0_s0_read;                // mm_interconnect_0:LCDFrameBuffer_0_s0_read -> LCDFrameBuffer_0:s0_read
	wire         mm_interconnect_0_lcdframebuffer_0_s0_write;               // mm_interconnect_0:LCDFrameBuffer_0_s0_write -> LCDFrameBuffer_0:s0_write
	wire  [31:0] mm_interconnect_0_lcdframebuffer_0_s0_writedata;           // mm_interconnect_0:LCDFrameBuffer_0_s0_writedata -> LCDFrameBuffer_0:s0_writedata
	wire         mm_interconnect_0_onchip_memory2_s1_chipselect;            // mm_interconnect_0:onchip_memory2_s1_chipselect -> onchip_memory2:chipselect
	wire  [31:0] mm_interconnect_0_onchip_memory2_s1_readdata;              // onchip_memory2:readdata -> mm_interconnect_0:onchip_memory2_s1_readdata
	wire  [15:0] mm_interconnect_0_onchip_memory2_s1_address;               // mm_interconnect_0:onchip_memory2_s1_address -> onchip_memory2:address
	wire   [3:0] mm_interconnect_0_onchip_memory2_s1_byteenable;            // mm_interconnect_0:onchip_memory2_s1_byteenable -> onchip_memory2:byteenable
	wire         mm_interconnect_0_onchip_memory2_s1_write;                 // mm_interconnect_0:onchip_memory2_s1_write -> onchip_memory2:write
	wire  [31:0] mm_interconnect_0_onchip_memory2_s1_writedata;             // mm_interconnect_0:onchip_memory2_s1_writedata -> onchip_memory2:writedata
	wire         mm_interconnect_0_onchip_memory2_s1_clken;                 // mm_interconnect_0:onchip_memory2_s1_clken -> onchip_memory2:clken
	wire         mm_interconnect_0_timer_0_s1_chipselect;                   // mm_interconnect_0:timer_0_s1_chipselect -> timer_0:chipselect
	wire  [15:0] mm_interconnect_0_timer_0_s1_readdata;                     // timer_0:readdata -> mm_interconnect_0:timer_0_s1_readdata
	wire   [2:0] mm_interconnect_0_timer_0_s1_address;                      // mm_interconnect_0:timer_0_s1_address -> timer_0:address
	wire         mm_interconnect_0_timer_0_s1_write;                        // mm_interconnect_0:timer_0_s1_write -> timer_0:write_n
	wire  [15:0] mm_interconnect_0_timer_0_s1_writedata;                    // mm_interconnect_0:timer_0_s1_writedata -> timer_0:writedata
	wire         mm_interconnect_0_spi_avalon_sd_0_sd_chipselect;           // mm_interconnect_0:SPI_AVALON_SD_0_sd_chipselect -> SPI_AVALON_SD_0:sd_chipselect
	wire  [31:0] mm_interconnect_0_spi_avalon_sd_0_sd_readdata;             // SPI_AVALON_SD_0:sd_readdata -> mm_interconnect_0:SPI_AVALON_SD_0_sd_readdata
	wire   [1:0] mm_interconnect_0_spi_avalon_sd_0_sd_address;              // mm_interconnect_0:SPI_AVALON_SD_0_sd_address -> SPI_AVALON_SD_0:sd_address
	wire         mm_interconnect_0_spi_avalon_sd_0_sd_write;                // mm_interconnect_0:SPI_AVALON_SD_0_sd_write -> SPI_AVALON_SD_0:sd_write
	wire  [31:0] mm_interconnect_0_spi_avalon_sd_0_sd_writedata;            // mm_interconnect_0:SPI_AVALON_SD_0_sd_writedata -> SPI_AVALON_SD_0:sd_writedata
	wire         irq_mapper_receiver0_irq;                                  // jtag_uart:av_irq -> irq_mapper:receiver0_irq
	wire  [31:0] cpu_irq_irq;                                               // irq_mapper:sender_irq -> cpu:irq
	wire         irq_mapper_receiver1_irq;                                  // irq_synchronizer:sender_irq -> irq_mapper:receiver1_irq
	wire   [0:0] irq_synchronizer_receiver_irq;                             // timer_0:irq -> irq_synchronizer:receiver_irq
	wire         irq_mapper_receiver2_irq;                                  // irq_synchronizer_001:sender_irq -> irq_mapper:receiver2_irq
	wire   [0:0] irq_synchronizer_001_receiver_irq;                         // dma_0:dma_ctl_irq -> irq_synchronizer_001:receiver_irq
	wire         rst_controller_reset_out_reset;                            // rst_controller:reset_out -> [LCDFrameBuffer_0:rst, dma_0:system_reset_n, irq_synchronizer:receiver_reset, irq_synchronizer_001:receiver_reset, mm_interconnect_0:LCDFrameBuffer_0_rst_reset_bridge_in_reset_reset, timer_0:reset_n]
	wire         rst_controller_001_reset_out_reset;                        // rst_controller_001:reset_out -> [SPI_AVALON_SD_0:reset, cpu:reset_n, i2c_AVALON_0:reset, irq_mapper:reset, irq_synchronizer:sender_reset, irq_synchronizer_001:sender_reset, jtag_uart:rst_n, mm_interconnect_0:cpu_reset_reset_bridge_in_reset_reset, new_sdram_controller_0:reset_n, onchip_memory2:reset, rst_translator:in_reset]
	wire         rst_controller_001_reset_out_reset_req;                    // rst_controller_001:reset_req -> [cpu:reset_req, onchip_memory2:reset_req, rst_translator:reset_req_in]

	LCD_AVALON lcdframebuffer_0 (
		.clk              (clk_clk),                                          //         clock.clk
		.s0_address       (mm_interconnect_0_lcdframebuffer_0_s0_address),    //            s0.address
		.s0_read          (mm_interconnect_0_lcdframebuffer_0_s0_read),       //              .read
		.s0_write         (mm_interconnect_0_lcdframebuffer_0_s0_write),      //              .write
		.s0_chipselect    (mm_interconnect_0_lcdframebuffer_0_s0_chipselect), //              .chipselect
		.s0_writedata     (mm_interconnect_0_lcdframebuffer_0_s0_writedata),  //              .writedata
		.s0_readdata      (mm_interconnect_0_lcdframebuffer_0_s0_readdata),   //              .readdata
		.lcd_cs           (lcd_lcd_cs),                                       //      External.lcd_cs
		.lcd_data         (lcd_lcd_data),                                     //              .lcd_data
		.lcd_dc           (lcd_lcd_dc),                                       //              .lcd_dc
		.lcd_rst          (lcd_lcd_rst),                                      //              .lcd_rst
		.lcd_wr           (lcd_lcd_wr),                                       //              .lcd_wr
		.rst              (rst_controller_reset_out_reset),                   //           rst.reset
		.m0_waitrequest   (lcdframebuffer_0_avalon_master_waitrequest),       // avalon_master.waitrequest
		.m0_readdatavalid (lcdframebuffer_0_avalon_master_readdatavalid),     //              .readdatavalid
		.m0_readdata      (lcdframebuffer_0_avalon_master_readdata),          //              .readdata
		.m0_address       (lcdframebuffer_0_avalon_master_address),           //              .address
		.m0_writedata     (lcdframebuffer_0_avalon_master_writedata),         //              .writedata
		.m0_chipselect    (lcdframebuffer_0_avalon_master_chipselect),        //              .chipselect
		.m0_byteenable_n  (lcdframebuffer_0_avalon_master_byteenable),        //              .byteenable_n
		.m0_read_n        (lcdframebuffer_0_avalon_master_read),              //              .read_n
		.m0_write_n       (lcdframebuffer_0_avalon_master_write)              //              .write_n
	);

	SPI_AVALON_SD spi_avalon_sd_0 (
		.clk           (pll_outclk0_clk),                                 //       clock.clk
		.reset         (rst_controller_001_reset_out_reset),              //       reset.reset
		.sd_chipselect (mm_interconnect_0_spi_avalon_sd_0_sd_chipselect), //          sd.chipselect
		.sd_write      (mm_interconnect_0_spi_avalon_sd_0_sd_write),      //            .write
		.sd_address    (mm_interconnect_0_spi_avalon_sd_0_sd_address),    //            .address
		.sd_writedata  (mm_interconnect_0_spi_avalon_sd_0_sd_writedata),  //            .writedata
		.sd_readdata   (mm_interconnect_0_spi_avalon_sd_0_sd_readdata),   //            .readdata
		.sd_cs         (sd_sd_cs),                                        // conduit_end.sd_cs
		.sd_clk        (sd_sd_clk),                                       //            .sd_clk
		.sd_di         (sd_sd_di),                                        //            .sd_di
		.sd_do         (sd_sd_do)                                         //            .sd_do
	);

	DE1_SOC_NIOS_2_cpu cpu (
		.clk                                 (pll_outclk0_clk),                                   //                       clk.clk
		.reset_n                             (~rst_controller_001_reset_out_reset),               //                     reset.reset_n
		.reset_req                           (rst_controller_001_reset_out_reset_req),            //                          .reset_req
		.d_address                           (cpu_data_master_address),                           //               data_master.address
		.d_byteenable                        (cpu_data_master_byteenable),                        //                          .byteenable
		.d_read                              (cpu_data_master_read),                              //                          .read
		.d_readdata                          (cpu_data_master_readdata),                          //                          .readdata
		.d_waitrequest                       (cpu_data_master_waitrequest),                       //                          .waitrequest
		.d_write                             (cpu_data_master_write),                             //                          .write
		.d_writedata                         (cpu_data_master_writedata),                         //                          .writedata
		.debug_mem_slave_debugaccess_to_roms (cpu_data_master_debugaccess),                       //                          .debugaccess
		.i_address                           (cpu_instruction_master_address),                    //        instruction_master.address
		.i_read                              (cpu_instruction_master_read),                       //                          .read
		.i_readdata                          (cpu_instruction_master_readdata),                   //                          .readdata
		.i_waitrequest                       (cpu_instruction_master_waitrequest),                //                          .waitrequest
		.irq                                 (cpu_irq_irq),                                       //                       irq.irq
		.debug_reset_request                 (),                                                  //       debug_reset_request.reset
		.debug_mem_slave_address             (mm_interconnect_0_cpu_debug_mem_slave_address),     //           debug_mem_slave.address
		.debug_mem_slave_byteenable          (mm_interconnect_0_cpu_debug_mem_slave_byteenable),  //                          .byteenable
		.debug_mem_slave_debugaccess         (mm_interconnect_0_cpu_debug_mem_slave_debugaccess), //                          .debugaccess
		.debug_mem_slave_read                (mm_interconnect_0_cpu_debug_mem_slave_read),        //                          .read
		.debug_mem_slave_readdata            (mm_interconnect_0_cpu_debug_mem_slave_readdata),    //                          .readdata
		.debug_mem_slave_waitrequest         (mm_interconnect_0_cpu_debug_mem_slave_waitrequest), //                          .waitrequest
		.debug_mem_slave_write               (mm_interconnect_0_cpu_debug_mem_slave_write),       //                          .write
		.debug_mem_slave_writedata           (mm_interconnect_0_cpu_debug_mem_slave_writedata),   //                          .writedata
		.dummy_ci_port                       ()                                                   // custom_instruction_master.readra
	);

	DE1_SOC_NIOS_2_dma_0 dma_0 (
		.clk                (clk_clk),                                               //                clk.clk
		.system_reset_n     (~rst_controller_reset_out_reset),                       //              reset.reset_n
		.dma_ctl_address    (mm_interconnect_0_dma_0_control_port_slave_address),    // control_port_slave.address
		.dma_ctl_chipselect (mm_interconnect_0_dma_0_control_port_slave_chipselect), //                   .chipselect
		.dma_ctl_readdata   (mm_interconnect_0_dma_0_control_port_slave_readdata),   //                   .readdata
		.dma_ctl_write_n    (~mm_interconnect_0_dma_0_control_port_slave_write),     //                   .write_n
		.dma_ctl_writedata  (mm_interconnect_0_dma_0_control_port_slave_writedata),  //                   .writedata
		.dma_ctl_irq        (irq_synchronizer_001_receiver_irq),                     //                irq.irq
		.read_address       (dma_0_read_master_address),                             //        read_master.address
		.read_chipselect    (dma_0_read_master_chipselect),                          //                   .chipselect
		.read_read_n        (dma_0_read_master_read),                                //                   .read_n
		.read_readdata      (dma_0_read_master_readdata),                            //                   .readdata
		.read_readdatavalid (dma_0_read_master_readdatavalid),                       //                   .readdatavalid
		.read_waitrequest   (dma_0_read_master_waitrequest),                         //                   .waitrequest
		.write_address      (dma_0_write_master_address),                            //       write_master.address
		.write_chipselect   (dma_0_write_master_chipselect),                         //                   .chipselect
		.write_waitrequest  (dma_0_write_master_waitrequest),                        //                   .waitrequest
		.write_write_n      (dma_0_write_master_write),                              //                   .write_n
		.write_writedata    (dma_0_write_master_writedata),                          //                   .writedata
		.write_byteenable   (dma_0_write_master_byteenable)                          //                   .byteenable
	);

	I2C_AVALON i2c_avalon_0 (
		.clk            (pll_outclk0_clk),                               //       clock.clk
		.reset          (rst_controller_001_reset_out_reset),            //       reset.reset
		.i2c_chipselect (mm_interconnect_0_i2c_avalon_0_i2c_chipselect), //         i2c.chipselect
		.i2c_write      (mm_interconnect_0_i2c_avalon_0_i2c_write),      //            .write
		.i2c_address    (mm_interconnect_0_i2c_avalon_0_i2c_address),    //            .address
		.i2c_writedata  (mm_interconnect_0_i2c_avalon_0_i2c_writedata),  //            .writedata
		.i2c_readdata   (mm_interconnect_0_i2c_avalon_0_i2c_readdata),   //            .readdata
		.i2c_reset      (i2c_rst),                                       // conduit_end.rst
		.i2c_sda        (i2c_sda),                                       //            .sda
		.i2c_sclk       (i2c_sclk)                                       //            .sclk
	);

	DE1_SOC_NIOS_2_jtag_uart jtag_uart (
		.clk            (pll_outclk0_clk),                                           //               clk.clk
		.rst_n          (~rst_controller_001_reset_out_reset),                       //             reset.reset_n
		.av_chipselect  (mm_interconnect_0_jtag_uart_avalon_jtag_slave_chipselect),  // avalon_jtag_slave.chipselect
		.av_address     (mm_interconnect_0_jtag_uart_avalon_jtag_slave_address),     //                  .address
		.av_read_n      (~mm_interconnect_0_jtag_uart_avalon_jtag_slave_read),       //                  .read_n
		.av_readdata    (mm_interconnect_0_jtag_uart_avalon_jtag_slave_readdata),    //                  .readdata
		.av_write_n     (~mm_interconnect_0_jtag_uart_avalon_jtag_slave_write),      //                  .write_n
		.av_writedata   (mm_interconnect_0_jtag_uart_avalon_jtag_slave_writedata),   //                  .writedata
		.av_waitrequest (mm_interconnect_0_jtag_uart_avalon_jtag_slave_waitrequest), //                  .waitrequest
		.av_irq         (irq_mapper_receiver0_irq)                                   //               irq.irq
	);

	DE1_SOC_NIOS_2_new_sdram_controller_0 new_sdram_controller_0 (
		.clk            (pll_outclk0_clk),                                           //   clk.clk
		.reset_n        (~rst_controller_001_reset_out_reset),                       // reset.reset_n
		.az_addr        (mm_interconnect_0_new_sdram_controller_0_s1_address),       //    s1.address
		.az_be_n        (~mm_interconnect_0_new_sdram_controller_0_s1_byteenable),   //      .byteenable_n
		.az_cs          (mm_interconnect_0_new_sdram_controller_0_s1_chipselect),    //      .chipselect
		.az_data        (mm_interconnect_0_new_sdram_controller_0_s1_writedata),     //      .writedata
		.az_rd_n        (~mm_interconnect_0_new_sdram_controller_0_s1_read),         //      .read_n
		.az_wr_n        (~mm_interconnect_0_new_sdram_controller_0_s1_write),        //      .write_n
		.za_data        (mm_interconnect_0_new_sdram_controller_0_s1_readdata),      //      .readdata
		.za_valid       (mm_interconnect_0_new_sdram_controller_0_s1_readdatavalid), //      .readdatavalid
		.za_waitrequest (mm_interconnect_0_new_sdram_controller_0_s1_waitrequest),   //      .waitrequest
		.zs_addr        (new_sdram_controller_0_wire_addr),                          //  wire.export
		.zs_ba          (new_sdram_controller_0_wire_ba),                            //      .export
		.zs_cas_n       (new_sdram_controller_0_wire_cas_n),                         //      .export
		.zs_cke         (new_sdram_controller_0_wire_cke),                           //      .export
		.zs_cs_n        (new_sdram_controller_0_wire_cs_n),                          //      .export
		.zs_dq          (new_sdram_controller_0_wire_dq),                            //      .export
		.zs_dqm         (new_sdram_controller_0_wire_dqm),                           //      .export
		.zs_ras_n       (new_sdram_controller_0_wire_ras_n),                         //      .export
		.zs_we_n        (new_sdram_controller_0_wire_we_n)                           //      .export
	);

	DE1_SOC_NIOS_2_onchip_memory2 onchip_memory2 (
		.clk        (pll_outclk0_clk),                                //   clk1.clk
		.address    (mm_interconnect_0_onchip_memory2_s1_address),    //     s1.address
		.clken      (mm_interconnect_0_onchip_memory2_s1_clken),      //       .clken
		.chipselect (mm_interconnect_0_onchip_memory2_s1_chipselect), //       .chipselect
		.write      (mm_interconnect_0_onchip_memory2_s1_write),      //       .write
		.readdata   (mm_interconnect_0_onchip_memory2_s1_readdata),   //       .readdata
		.writedata  (mm_interconnect_0_onchip_memory2_s1_writedata),  //       .writedata
		.byteenable (mm_interconnect_0_onchip_memory2_s1_byteenable), //       .byteenable
		.reset      (rst_controller_001_reset_out_reset),             // reset1.reset
		.reset_req  (rst_controller_001_reset_out_reset_req)          //       .reset_req
	);

	DE1_SOC_NIOS_2_pll pll (
		.refclk   (clk_clk),         //  refclk.clk
		.rst      (~reset_reset_n),  //   reset.reset
		.outclk_0 (pll_outclk0_clk), // outclk0.clk
		.outclk_1 (sdram_clk_clk),   // outclk1.clk
		.locked   ()                 // (terminated)
	);

	DE1_SOC_NIOS_2_timer_0 timer_0 (
		.clk        (clk_clk),                                 //   clk.clk
		.reset_n    (~rst_controller_reset_out_reset),         // reset.reset_n
		.address    (mm_interconnect_0_timer_0_s1_address),    //    s1.address
		.writedata  (mm_interconnect_0_timer_0_s1_writedata),  //      .writedata
		.readdata   (mm_interconnect_0_timer_0_s1_readdata),   //      .readdata
		.chipselect (mm_interconnect_0_timer_0_s1_chipselect), //      .chipselect
		.write_n    (~mm_interconnect_0_timer_0_s1_write),     //      .write_n
		.irq        (irq_synchronizer_receiver_irq)            //   irq.irq
	);

	DE1_SOC_NIOS_2_mm_interconnect_0 mm_interconnect_0 (
		.clk_0_clk_clk                                    (clk_clk),                                                   //                                  clk_0_clk.clk
		.pll_outclk0_clk                                  (pll_outclk0_clk),                                           //                                pll_outclk0.clk
		.cpu_reset_reset_bridge_in_reset_reset            (rst_controller_001_reset_out_reset),                        //            cpu_reset_reset_bridge_in_reset.reset
		.LCDFrameBuffer_0_rst_reset_bridge_in_reset_reset (rst_controller_reset_out_reset),                            // LCDFrameBuffer_0_rst_reset_bridge_in_reset.reset
		.cpu_data_master_address                          (cpu_data_master_address),                                   //                            cpu_data_master.address
		.cpu_data_master_waitrequest                      (cpu_data_master_waitrequest),                               //                                           .waitrequest
		.cpu_data_master_byteenable                       (cpu_data_master_byteenable),                                //                                           .byteenable
		.cpu_data_master_read                             (cpu_data_master_read),                                      //                                           .read
		.cpu_data_master_readdata                         (cpu_data_master_readdata),                                  //                                           .readdata
		.cpu_data_master_write                            (cpu_data_master_write),                                     //                                           .write
		.cpu_data_master_writedata                        (cpu_data_master_writedata),                                 //                                           .writedata
		.cpu_data_master_debugaccess                      (cpu_data_master_debugaccess),                               //                                           .debugaccess
		.cpu_instruction_master_address                   (cpu_instruction_master_address),                            //                     cpu_instruction_master.address
		.cpu_instruction_master_waitrequest               (cpu_instruction_master_waitrequest),                        //                                           .waitrequest
		.cpu_instruction_master_read                      (cpu_instruction_master_read),                               //                                           .read
		.cpu_instruction_master_readdata                  (cpu_instruction_master_readdata),                           //                                           .readdata
		.dma_0_read_master_address                        (dma_0_read_master_address),                                 //                          dma_0_read_master.address
		.dma_0_read_master_waitrequest                    (dma_0_read_master_waitrequest),                             //                                           .waitrequest
		.dma_0_read_master_chipselect                     (dma_0_read_master_chipselect),                              //                                           .chipselect
		.dma_0_read_master_read                           (~dma_0_read_master_read),                                   //                                           .read
		.dma_0_read_master_readdata                       (dma_0_read_master_readdata),                                //                                           .readdata
		.dma_0_read_master_readdatavalid                  (dma_0_read_master_readdatavalid),                           //                                           .readdatavalid
		.dma_0_write_master_address                       (dma_0_write_master_address),                                //                         dma_0_write_master.address
		.dma_0_write_master_waitrequest                   (dma_0_write_master_waitrequest),                            //                                           .waitrequest
		.dma_0_write_master_byteenable                    (dma_0_write_master_byteenable),                             //                                           .byteenable
		.dma_0_write_master_chipselect                    (dma_0_write_master_chipselect),                             //                                           .chipselect
		.dma_0_write_master_write                         (~dma_0_write_master_write),                                 //                                           .write
		.dma_0_write_master_writedata                     (dma_0_write_master_writedata),                              //                                           .writedata
		.LCDFrameBuffer_0_avalon_master_address           (lcdframebuffer_0_avalon_master_address),                    //             LCDFrameBuffer_0_avalon_master.address
		.LCDFrameBuffer_0_avalon_master_waitrequest       (lcdframebuffer_0_avalon_master_waitrequest),                //                                           .waitrequest
		.LCDFrameBuffer_0_avalon_master_byteenable        (~lcdframebuffer_0_avalon_master_byteenable),                //                                           .byteenable
		.LCDFrameBuffer_0_avalon_master_chipselect        (lcdframebuffer_0_avalon_master_chipselect),                 //                                           .chipselect
		.LCDFrameBuffer_0_avalon_master_read              (~lcdframebuffer_0_avalon_master_read),                      //                                           .read
		.LCDFrameBuffer_0_avalon_master_readdata          (lcdframebuffer_0_avalon_master_readdata),                   //                                           .readdata
		.LCDFrameBuffer_0_avalon_master_readdatavalid     (lcdframebuffer_0_avalon_master_readdatavalid),              //                                           .readdatavalid
		.LCDFrameBuffer_0_avalon_master_write             (~lcdframebuffer_0_avalon_master_write),                     //                                           .write
		.LCDFrameBuffer_0_avalon_master_writedata         (lcdframebuffer_0_avalon_master_writedata),                  //                                           .writedata
		.cpu_debug_mem_slave_address                      (mm_interconnect_0_cpu_debug_mem_slave_address),             //                        cpu_debug_mem_slave.address
		.cpu_debug_mem_slave_write                        (mm_interconnect_0_cpu_debug_mem_slave_write),               //                                           .write
		.cpu_debug_mem_slave_read                         (mm_interconnect_0_cpu_debug_mem_slave_read),                //                                           .read
		.cpu_debug_mem_slave_readdata                     (mm_interconnect_0_cpu_debug_mem_slave_readdata),            //                                           .readdata
		.cpu_debug_mem_slave_writedata                    (mm_interconnect_0_cpu_debug_mem_slave_writedata),           //                                           .writedata
		.cpu_debug_mem_slave_byteenable                   (mm_interconnect_0_cpu_debug_mem_slave_byteenable),          //                                           .byteenable
		.cpu_debug_mem_slave_waitrequest                  (mm_interconnect_0_cpu_debug_mem_slave_waitrequest),         //                                           .waitrequest
		.cpu_debug_mem_slave_debugaccess                  (mm_interconnect_0_cpu_debug_mem_slave_debugaccess),         //                                           .debugaccess
		.dma_0_control_port_slave_address                 (mm_interconnect_0_dma_0_control_port_slave_address),        //                   dma_0_control_port_slave.address
		.dma_0_control_port_slave_write                   (mm_interconnect_0_dma_0_control_port_slave_write),          //                                           .write
		.dma_0_control_port_slave_readdata                (mm_interconnect_0_dma_0_control_port_slave_readdata),       //                                           .readdata
		.dma_0_control_port_slave_writedata               (mm_interconnect_0_dma_0_control_port_slave_writedata),      //                                           .writedata
		.dma_0_control_port_slave_chipselect              (mm_interconnect_0_dma_0_control_port_slave_chipselect),     //                                           .chipselect
		.i2c_AVALON_0_i2c_address                         (mm_interconnect_0_i2c_avalon_0_i2c_address),                //                           i2c_AVALON_0_i2c.address
		.i2c_AVALON_0_i2c_write                           (mm_interconnect_0_i2c_avalon_0_i2c_write),                  //                                           .write
		.i2c_AVALON_0_i2c_readdata                        (mm_interconnect_0_i2c_avalon_0_i2c_readdata),               //                                           .readdata
		.i2c_AVALON_0_i2c_writedata                       (mm_interconnect_0_i2c_avalon_0_i2c_writedata),              //                                           .writedata
		.i2c_AVALON_0_i2c_chipselect                      (mm_interconnect_0_i2c_avalon_0_i2c_chipselect),             //                                           .chipselect
		.jtag_uart_avalon_jtag_slave_address              (mm_interconnect_0_jtag_uart_avalon_jtag_slave_address),     //                jtag_uart_avalon_jtag_slave.address
		.jtag_uart_avalon_jtag_slave_write                (mm_interconnect_0_jtag_uart_avalon_jtag_slave_write),       //                                           .write
		.jtag_uart_avalon_jtag_slave_read                 (mm_interconnect_0_jtag_uart_avalon_jtag_slave_read),        //                                           .read
		.jtag_uart_avalon_jtag_slave_readdata             (mm_interconnect_0_jtag_uart_avalon_jtag_slave_readdata),    //                                           .readdata
		.jtag_uart_avalon_jtag_slave_writedata            (mm_interconnect_0_jtag_uart_avalon_jtag_slave_writedata),   //                                           .writedata
		.jtag_uart_avalon_jtag_slave_waitrequest          (mm_interconnect_0_jtag_uart_avalon_jtag_slave_waitrequest), //                                           .waitrequest
		.jtag_uart_avalon_jtag_slave_chipselect           (mm_interconnect_0_jtag_uart_avalon_jtag_slave_chipselect),  //                                           .chipselect
		.LCDFrameBuffer_0_s0_address                      (mm_interconnect_0_lcdframebuffer_0_s0_address),             //                        LCDFrameBuffer_0_s0.address
		.LCDFrameBuffer_0_s0_write                        (mm_interconnect_0_lcdframebuffer_0_s0_write),               //                                           .write
		.LCDFrameBuffer_0_s0_read                         (mm_interconnect_0_lcdframebuffer_0_s0_read),                //                                           .read
		.LCDFrameBuffer_0_s0_readdata                     (mm_interconnect_0_lcdframebuffer_0_s0_readdata),            //                                           .readdata
		.LCDFrameBuffer_0_s0_writedata                    (mm_interconnect_0_lcdframebuffer_0_s0_writedata),           //                                           .writedata
		.LCDFrameBuffer_0_s0_chipselect                   (mm_interconnect_0_lcdframebuffer_0_s0_chipselect),          //                                           .chipselect
		.new_sdram_controller_0_s1_address                (mm_interconnect_0_new_sdram_controller_0_s1_address),       //                  new_sdram_controller_0_s1.address
		.new_sdram_controller_0_s1_write                  (mm_interconnect_0_new_sdram_controller_0_s1_write),         //                                           .write
		.new_sdram_controller_0_s1_read                   (mm_interconnect_0_new_sdram_controller_0_s1_read),          //                                           .read
		.new_sdram_controller_0_s1_readdata               (mm_interconnect_0_new_sdram_controller_0_s1_readdata),      //                                           .readdata
		.new_sdram_controller_0_s1_writedata              (mm_interconnect_0_new_sdram_controller_0_s1_writedata),     //                                           .writedata
		.new_sdram_controller_0_s1_byteenable             (mm_interconnect_0_new_sdram_controller_0_s1_byteenable),    //                                           .byteenable
		.new_sdram_controller_0_s1_readdatavalid          (mm_interconnect_0_new_sdram_controller_0_s1_readdatavalid), //                                           .readdatavalid
		.new_sdram_controller_0_s1_waitrequest            (mm_interconnect_0_new_sdram_controller_0_s1_waitrequest),   //                                           .waitrequest
		.new_sdram_controller_0_s1_chipselect             (mm_interconnect_0_new_sdram_controller_0_s1_chipselect),    //                                           .chipselect
		.onchip_memory2_s1_address                        (mm_interconnect_0_onchip_memory2_s1_address),               //                          onchip_memory2_s1.address
		.onchip_memory2_s1_write                          (mm_interconnect_0_onchip_memory2_s1_write),                 //                                           .write
		.onchip_memory2_s1_readdata                       (mm_interconnect_0_onchip_memory2_s1_readdata),              //                                           .readdata
		.onchip_memory2_s1_writedata                      (mm_interconnect_0_onchip_memory2_s1_writedata),             //                                           .writedata
		.onchip_memory2_s1_byteenable                     (mm_interconnect_0_onchip_memory2_s1_byteenable),            //                                           .byteenable
		.onchip_memory2_s1_chipselect                     (mm_interconnect_0_onchip_memory2_s1_chipselect),            //                                           .chipselect
		.onchip_memory2_s1_clken                          (mm_interconnect_0_onchip_memory2_s1_clken),                 //                                           .clken
		.SPI_AVALON_SD_0_sd_address                       (mm_interconnect_0_spi_avalon_sd_0_sd_address),              //                         SPI_AVALON_SD_0_sd.address
		.SPI_AVALON_SD_0_sd_write                         (mm_interconnect_0_spi_avalon_sd_0_sd_write),                //                                           .write
		.SPI_AVALON_SD_0_sd_readdata                      (mm_interconnect_0_spi_avalon_sd_0_sd_readdata),             //                                           .readdata
		.SPI_AVALON_SD_0_sd_writedata                     (mm_interconnect_0_spi_avalon_sd_0_sd_writedata),            //                                           .writedata
		.SPI_AVALON_SD_0_sd_chipselect                    (mm_interconnect_0_spi_avalon_sd_0_sd_chipselect),           //                                           .chipselect
		.timer_0_s1_address                               (mm_interconnect_0_timer_0_s1_address),                      //                                 timer_0_s1.address
		.timer_0_s1_write                                 (mm_interconnect_0_timer_0_s1_write),                        //                                           .write
		.timer_0_s1_readdata                              (mm_interconnect_0_timer_0_s1_readdata),                     //                                           .readdata
		.timer_0_s1_writedata                             (mm_interconnect_0_timer_0_s1_writedata),                    //                                           .writedata
		.timer_0_s1_chipselect                            (mm_interconnect_0_timer_0_s1_chipselect)                    //                                           .chipselect
	);

	DE1_SOC_NIOS_2_irq_mapper irq_mapper (
		.clk           (pll_outclk0_clk),                    //       clk.clk
		.reset         (rst_controller_001_reset_out_reset), // clk_reset.reset
		.receiver0_irq (irq_mapper_receiver0_irq),           // receiver0.irq
		.receiver1_irq (irq_mapper_receiver1_irq),           // receiver1.irq
		.receiver2_irq (irq_mapper_receiver2_irq),           // receiver2.irq
		.sender_irq    (cpu_irq_irq)                         //    sender.irq
	);

	altera_irq_clock_crosser #(
		.IRQ_WIDTH (1)
	) irq_synchronizer (
		.receiver_clk   (clk_clk),                            //       receiver_clk.clk
		.sender_clk     (pll_outclk0_clk),                    //         sender_clk.clk
		.receiver_reset (rst_controller_reset_out_reset),     // receiver_clk_reset.reset
		.sender_reset   (rst_controller_001_reset_out_reset), //   sender_clk_reset.reset
		.receiver_irq   (irq_synchronizer_receiver_irq),      //           receiver.irq
		.sender_irq     (irq_mapper_receiver1_irq)            //             sender.irq
	);

	altera_irq_clock_crosser #(
		.IRQ_WIDTH (1)
	) irq_synchronizer_001 (
		.receiver_clk   (clk_clk),                            //       receiver_clk.clk
		.sender_clk     (pll_outclk0_clk),                    //         sender_clk.clk
		.receiver_reset (rst_controller_reset_out_reset),     // receiver_clk_reset.reset
		.sender_reset   (rst_controller_001_reset_out_reset), //   sender_clk_reset.reset
		.receiver_irq   (irq_synchronizer_001_receiver_irq),  //           receiver.irq
		.sender_irq     (irq_mapper_receiver2_irq)            //             sender.irq
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller (
		.reset_in0      (~reset_reset_n),                 // reset_in0.reset
		.clk            (clk_clk),                        //       clk.clk
		.reset_out      (rst_controller_reset_out_reset), // reset_out.reset
		.reset_req      (),                               // (terminated)
		.reset_req_in0  (1'b0),                           // (terminated)
		.reset_in1      (1'b0),                           // (terminated)
		.reset_req_in1  (1'b0),                           // (terminated)
		.reset_in2      (1'b0),                           // (terminated)
		.reset_req_in2  (1'b0),                           // (terminated)
		.reset_in3      (1'b0),                           // (terminated)
		.reset_req_in3  (1'b0),                           // (terminated)
		.reset_in4      (1'b0),                           // (terminated)
		.reset_req_in4  (1'b0),                           // (terminated)
		.reset_in5      (1'b0),                           // (terminated)
		.reset_req_in5  (1'b0),                           // (terminated)
		.reset_in6      (1'b0),                           // (terminated)
		.reset_req_in6  (1'b0),                           // (terminated)
		.reset_in7      (1'b0),                           // (terminated)
		.reset_req_in7  (1'b0),                           // (terminated)
		.reset_in8      (1'b0),                           // (terminated)
		.reset_req_in8  (1'b0),                           // (terminated)
		.reset_in9      (1'b0),                           // (terminated)
		.reset_req_in9  (1'b0),                           // (terminated)
		.reset_in10     (1'b0),                           // (terminated)
		.reset_req_in10 (1'b0),                           // (terminated)
		.reset_in11     (1'b0),                           // (terminated)
		.reset_req_in11 (1'b0),                           // (terminated)
		.reset_in12     (1'b0),                           // (terminated)
		.reset_req_in12 (1'b0),                           // (terminated)
		.reset_in13     (1'b0),                           // (terminated)
		.reset_req_in13 (1'b0),                           // (terminated)
		.reset_in14     (1'b0),                           // (terminated)
		.reset_req_in14 (1'b0),                           // (terminated)
		.reset_in15     (1'b0),                           // (terminated)
		.reset_req_in15 (1'b0)                            // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (1),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_001 (
		.reset_in0      (~reset_reset_n),                         // reset_in0.reset
		.clk            (pll_outclk0_clk),                        //       clk.clk
		.reset_out      (rst_controller_001_reset_out_reset),     // reset_out.reset
		.reset_req      (rst_controller_001_reset_out_reset_req), //          .reset_req
		.reset_req_in0  (1'b0),                                   // (terminated)
		.reset_in1      (1'b0),                                   // (terminated)
		.reset_req_in1  (1'b0),                                   // (terminated)
		.reset_in2      (1'b0),                                   // (terminated)
		.reset_req_in2  (1'b0),                                   // (terminated)
		.reset_in3      (1'b0),                                   // (terminated)
		.reset_req_in3  (1'b0),                                   // (terminated)
		.reset_in4      (1'b0),                                   // (terminated)
		.reset_req_in4  (1'b0),                                   // (terminated)
		.reset_in5      (1'b0),                                   // (terminated)
		.reset_req_in5  (1'b0),                                   // (terminated)
		.reset_in6      (1'b0),                                   // (terminated)
		.reset_req_in6  (1'b0),                                   // (terminated)
		.reset_in7      (1'b0),                                   // (terminated)
		.reset_req_in7  (1'b0),                                   // (terminated)
		.reset_in8      (1'b0),                                   // (terminated)
		.reset_req_in8  (1'b0),                                   // (terminated)
		.reset_in9      (1'b0),                                   // (terminated)
		.reset_req_in9  (1'b0),                                   // (terminated)
		.reset_in10     (1'b0),                                   // (terminated)
		.reset_req_in10 (1'b0),                                   // (terminated)
		.reset_in11     (1'b0),                                   // (terminated)
		.reset_req_in11 (1'b0),                                   // (terminated)
		.reset_in12     (1'b0),                                   // (terminated)
		.reset_req_in12 (1'b0),                                   // (terminated)
		.reset_in13     (1'b0),                                   // (terminated)
		.reset_req_in13 (1'b0),                                   // (terminated)
		.reset_in14     (1'b0),                                   // (terminated)
		.reset_req_in14 (1'b0),                                   // (terminated)
		.reset_in15     (1'b0),                                   // (terminated)
		.reset_req_in15 (1'b0)                                    // (terminated)
	);

endmodule
